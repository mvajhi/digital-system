module ShiftReg (
    input wire clk,
    input wire reset,
    input wire load,
    input wire shift_in,
    output wire [15:0] shift_out
);

    reg [15:0] reg;

    always @(posedge clk or posedge reset) begin
        if (reset)
            reg <= 16'b0;
        else if (load)
            reg <= shift_in;
        else
            reg <= {reg[14:0], 1'b0};
    end

    assign shift_out = reg;

endmodule